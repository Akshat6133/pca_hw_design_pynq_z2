
module fifo (
    input  wire clk,
    input  wire rst_n
);
    // Placeholder – real logic later
endmodule
